imperative-edsl-vhdl
