york-lava
