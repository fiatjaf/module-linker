clash-vhdl
